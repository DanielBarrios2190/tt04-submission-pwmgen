`timescale 1ns / 1ps

module tt_um_db_PWM(
    input  wire [7:0] ui_in,    // Dedicated inputs - connected to the input switches
    output wire [7:0] uo_out,   // Dedicated outputs - connected to the 7 segment display
    input  wire [7:0] uio_in,   // IOs: Bidirectional Input path
    output wire [7:0] uio_out,  // IOs: Bidirectional Output path
    output wire [7:0] uio_oe,   // IOs: Bidirectional Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // will go high when the design is enabled
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset

    );
    parameter BITS_duty = 3;
    wire clk_in;
    wire rst;
    wire [BITS_duty:0] duty;
    //wire pwm_out;

    assign duty = ui_in[BITS_duty:0];
    assign clk_in = clk;
    assign rst = ~rst_n;

    reg [BITS_duty:0] cnt;
    //reg pwm_q;
    //wire pwm_d;

    //assign pwm_d = (cnt < duty);  
    
    always @(posedge clk_in or posedge rst) begin
        if(rst) begin
         //pwm_q <=0;
         cnt <= 0;
        end else begin
         //pwm_q <= pwm_d;
         
         if((cnt >= (2**BITS_duty)-1))
            cnt <= 0;
         else begin      
            cnt <= cnt + 1;
         end
        end
    end

    assign uo_out[0] = (cnt < duty);

endmodule
